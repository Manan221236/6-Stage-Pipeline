// SYNCHRONIZED TESTBENCH for 6-Stage Pipeline K²RED Implementation
// Perfectly aligned with instruction memory layout

module K2RED_Dilithium_tb;

    //---------------------------- 1. Clock & Reset ----------------------------
    reg  clk;
    reg  rst;                     // active-HIGH reset
    
    initial begin
        clk = 0;
        forever #10 clk = ~clk;   // 50 MHz clock
    end
    
    //---------------------------- 2. Debug Signal Wires -----------------------
    wire [31:0] debug_alu_result;
    wire [4:0]  debug_reg_addr;
    wire        debug_reg_write;
    wire        debug_mem_write;

    //---------------------------- 3. Device Under Test ------------------------
    Pipeline_top dut ( 
        .clk(clk), 
        .rst(rst),
        .debug_alu_result(debug_alu_result),
        .debug_reg_addr(debug_reg_addr),
        .debug_reg_write(debug_reg_write),
        .debug_mem_write(debug_mem_write)
    );

    //---------------------------- 4. Simulation Setup -------------------------
    initial begin
        $dumpfile("k2red_dilithium_6stage.vcd");
        $dumpvars(0, K2RED_Dilithium_tb);
        
        // Explicitly dump debug signals
        $dumpvars(1, debug_alu_result, debug_reg_addr, debug_reg_write, debug_mem_write);
        
        // Reset sequence
        rst = 1;  
        repeat (5) @(posedge clk);   // 5 cycles reset
        rst = 0;                     // release reset
        
        $display("=== K²RED CRYSTALS-DILITHIUM TEST (6-STAGE SYNCHRONIZED) ===");
        $display("Testing: K²RED modular multiplication with Dilithium parameters");
        $display("Parameters: P=8380417, k=1023, m=13, n=24");
        $display("Pipeline: 6-stage with synchronized NOP timing");
        $display("Input: A=12345, B=6789, Expected A*B=83810205");
        $display("Termination: ECALL at address 0xA0 (mem[64])");
    end

    //---------------------------- 5. Cycle Counter ----------------------------
    integer cyc;
    initial cyc = 0;
    always @(posedge clk) begin
        if (!rst) cyc = cyc + 1;
    end

    //---------------------------- 6. Basic Debug Output -----------------------
    always @(posedge clk) begin
        if (!rst) begin
            $display("DEBUG: cyc=%0d alu_result=0x%08h reg_addr=x%0d reg_write=%b mem_write=%b",
                     cyc, debug_alu_result, debug_reg_addr, debug_reg_write, debug_mem_write);
        end
    end

    //---------------------------- 7. Register Monitoring ----------------------
    always @(posedge clk) begin
        if (!rst && (cyc % 25 == 0) && (cyc > 0)) begin  // Every 25 cycles
            $display("DILITHIUM_REGS: cyc=%0d x10=%0d x12=%0d x14=%0d x15=%0d x16=%0d x24=%0d x7=%0d", 
                     cyc, $signed(dut.Decode.rf.regf[10]), $signed(dut.Decode.rf.regf[12]),
                     $signed(dut.Decode.rf.regf[14]), $signed(dut.Decode.rf.regf[15]),
                     $signed(dut.Decode.rf.regf[16]), $signed(dut.Decode.rf.regf[24]), 
                     $signed(dut.Decode.rf.regf[7]));
        end
    end

    //---------------------------- 8. SYNCHRONIZED Phase Detection (UPDATED) ---
    reg [3:0] test_phase;
    initial test_phase = 0;
    
    always @(posedge clk) begin
        if (!rst) begin
            case (dut.PCD)
                // UPDATED: Synchronized with new instruction memory layout
                32'h00000000: test_phase = 1;  // Phase 1: Parameter setup (0x00-0x24)
                32'h00000028: test_phase = 2;  // Phase 2: Input values (0x28-0x54) - EXTENDED
                32'h00000058: test_phase = 3;  // Phase 3: K²RED algorithm (0x58-0xF0) - SHIFTED
                32'h000000F4: test_phase = 4;  // Phase 4: Test validation (0xF4-0x108) - SHIFTED
                32'h00000110: test_phase = 5;  // Phase 5: Program termination (0x110) - SHIFTED
            endcase
        end
    end
    
    // Phase change detection
    reg [3:0] prev_test_phase;
    always @(posedge clk) begin
        if (!rst) begin
            if (test_phase != prev_test_phase) begin
                case (test_phase)
                    1: $display("\n=== PHASE 1: PARAMETER SETUP (0x00-0x24) ===");
                    2: $display("\n=== PHASE 2: INPUT VALUES (0x28-0x54) EXTENDED ===");
                    3: $display("\n=== PHASE 3: K²RED ALGORITHM (0x58-0xF0) SHIFTED ===");
                    4: $display("\n=== PHASE 4: TEST VALIDATION (0xF4-0x108) SHIFTED ===");
                    5: $display("\n=== PHASE 5: PROGRAM TERMINATION (0x110) SHIFTED ===");
                endcase
                prev_test_phase = test_phase;
            end
        end
    end

    //---------------------------- 9. Value Validation -------------------------
    always @(posedge clk) begin
        if (!rst && debug_reg_write && (debug_reg_addr != 5'd0)) begin
            case (debug_reg_addr)
                // Parameters
                5'd10: begin
                    $display("DILITHIUM: k <= %0d (parameter k=1023)", $signed(debug_alu_result));
                    if (debug_alu_result == 32'd1023) 
                        $display("✅ CORRECT: k=1023 loaded successfully");
                end
                5'd11: begin
                    $display("DILITHIUM: m <= %0d (parameter m=13)", $signed(debug_alu_result));
                    if (debug_alu_result == 32'd13) 
                        $display("✅ CORRECT: m=13 loaded successfully");
                end
                5'd12: begin
                    $display("DILITHIUM: P <= %0d (parameter P=8380417)", $signed(debug_alu_result));
                    if (debug_alu_result == 32'd8380417) 
                        $display("✅ CORRECT: P=8380417 loaded successfully");
                end
                5'd13: begin
                    $display("DILITHIUM: n <= %0d (parameter n=24)", $signed(debug_alu_result));
                    if (debug_alu_result == 32'd24) 
                        $display("✅ CORRECT: n=24 loaded successfully");
                end
                
                // Input values - CRITICAL VALIDATION
                5'd14: begin
                    $display("DILITHIUM: A <= %0d (input A=12345)", $signed(debug_alu_result));
                    if (debug_alu_result == 32'd12345) 
                        $display("✅ PERFECT: A=12345 loaded correctly!");
                    else 
                        $display("❌ ERROR: A=%0d, expected 12345", $signed(debug_alu_result));
                end
                5'd15: begin
                    $display("DILITHIUM: B <= %0d (input B=6789)", $signed(debug_alu_result));
                    if (debug_alu_result == 32'd6789) 
                        $display("✅ PERFECT: B=6789 loaded correctly!");
                    else 
                        $display("❌ ERROR: B=%0d, expected 6789", $signed(debug_alu_result));
                end
                
                // Computation results
                5'd16: begin
                    $display("DILITHIUM: R_low <= %0d (A*B lower 32 bits)", $signed(debug_alu_result));
                    if (debug_alu_result == 32'd83810205) 
                        $display("✅ PERFECT: A*B=83810205 (12345*6789) correct!");
                    else 
                        $display("❌ ERROR: A*B=%0d, expected 83810205", $signed(debug_alu_result));
                end
                5'd17: $display("DILITHIUM: R_high <= %0d (A*B upper 32 bits)", $signed(debug_alu_result));
                5'd18: $display("DILITHIUM: Rl <= %0d (lower 13 bits)", $signed(debug_alu_result));
                5'd19: $display("DILITHIUM: Rh <= %0d (upper bits)", $signed(debug_alu_result));
                5'd20: $display("DILITHIUM: C <= %0d (k*Rl - Rh)", $signed(debug_alu_result));
                5'd21: $display("DILITHIUM: Cl <= %0d (lower 13 bits of C)", $signed(debug_alu_result));
                5'd22: $display("DILITHIUM: Ch <= %0d (upper bits of C)", $signed(debug_alu_result));
                5'd23: $display("DILITHIUM: C' <= %0d (INTERMEDIATE RESULT)", $signed(debug_alu_result));
                5'd24: begin
                    $display("DILITHIUM: FINAL RESULT <= %0d (0x%08h)", $signed(debug_alu_result), debug_alu_result);
                    if (debug_alu_result != 32'd0) 
                        $display("✅ SUCCESS: K²RED algorithm produced non-zero result!");
                    else 
                        $display("❌ WARNING: K²RED result is zero");
                end
                
                // Test validation
                5'd7: begin
                    $display("VALIDATION: Test counter <= %0d (should reach 5)", $signed(debug_alu_result));
                    if (debug_alu_result == 32'd5) 
                        $display("✅ SUCCESS: Test counter reached 5!");
                    else if (debug_alu_result > 0) 
                        $display("🔄 PROGRESS: Test counter = %0d", $signed(debug_alu_result));
                end
                
                default: $display("REGWRITE: x%0d <= %0d (0x%08h)", 
                                debug_reg_addr, $signed(debug_alu_result), debug_alu_result);
            endcase
        end
    end

    //---------------------------- 10. Multiplication Detection ----------------
    always @(posedge clk) begin
        if (!rst && (dut.InstrD[6:0] == 7'b0110011) && (dut.InstrD[31:25] == 7'b0000001)) begin
            case (dut.InstrD[14:12])
                3'b000: $display("DILITHIUM_MUL: MUL instruction at PC=0x%08h", dut.PCD);
                3'b001: $display("DILITHIUM_MULH: MULH instruction at PC=0x%08h", dut.PCD);
            endcase
        end
    end

    //---------------------------- 11. Instruction Trace -----------------------
    integer trace_log;
    initial begin
        trace_log = $fopen("k2red_dilithium_sync_trace.txt", "w");
    end
    
    always @(posedge clk) begin
        if (!rst && (dut.InstrD != 32'h0000_0013)) begin
            $display("TRACE: cyc=%0d PC=0x%08h instr=0x%08h", cyc, dut.PCD, dut.InstrD);
            $fdisplay(trace_log, "%0d,0x%08h,0x%08h", cyc, dut.PCD, dut.InstrD);
        end
    end

    //---------------------------- 12. Comprehensive Result Verification -------
    task verify_dilithium_results;
        reg [31:0] k2red_result, test_counter;
        reg [31:0] k_param, p_param, m_param, n_param;
        reg [31:0] input_a, input_b, mult_result_low, mult_result_high;
        integer errors, warnings;
        begin
            // Read all critical registers
            k2red_result = dut.Decode.rf.regf[24];      // Final K²RED result
            test_counter = dut.Decode.rf.regf[7];       // Test validation counter
            k_param = dut.Decode.rf.regf[10];           // k parameter
            p_param = dut.Decode.rf.regf[12];           // P parameter  
            m_param = dut.Decode.rf.regf[11];           // m parameter
            n_param = dut.Decode.rf.regf[13];           // n parameter
            input_a = dut.Decode.rf.regf[14];           // Input A
            input_b = dut.Decode.rf.regf[15];           // Input B
            mult_result_low = dut.Decode.rf.regf[16];   // A*B lower 32 bits
            mult_result_high = dut.Decode.rf.regf[17];  // A*B upper 32 bits
            
            errors = 0;
            warnings = 0;
            
            $display("\n" + "="*80);
            $display("K²RED CRYSTALS-DILITHIUM SYNCHRONIZED TEST RESULTS");
            $display("="*80);
            
            $display("\n📊 ALGORITHM PARAMETERS:");
            $display("  k = %0d (expected: 1023)", k_param);
            $display("  P = %0d (expected: 8380417)", p_param);
            $display("  m = %0d (expected: 13)", m_param);
            $display("  n = %0d (expected: 24)", n_param);
            
            $display("\n🔢 INPUT VALUES:");
            $display("  A = %0d (expected: 12345)", $signed(input_a));
            $display("  B = %0d (expected: 6789)", $signed(input_b));
            
            $display("\n🧮 COMPUTATION RESULTS:");
            $display("  A*B (low)  = %0d (expected: 83810205)", $signed(mult_result_low));
            $display("  A*B (high) = %0d (expected: 0)", $signed(mult_result_high));
            $display("  K²RED      = %0d (0x%08h)", $signed(k2red_result), k2red_result);
            $display("  Test count = %0d (expected: 5)", test_counter);
            
            $display("\n🔍 DETAILED VALIDATION:");
            
            // Parameter validation
            if (k_param !== 32'd1023) begin
                $display("❌ FAIL: k parameter incorrect");
                errors = errors + 1;
            end else $display("✅ PASS: k=1023 parameter correct");
            
            if (p_param !== 32'd8380417) begin
                $display("❌ FAIL: P parameter incorrect");
                errors = errors + 1;
            end else $display("✅ PASS: P=8380417 parameter correct");
            
            if (m_param !== 32'd13) begin
                $display("❌ FAIL: m parameter incorrect");
                errors = errors + 1;
            end else $display("✅ PASS: m=13 parameter correct");
            
            if (n_param !== 32'd24) begin
                $display("❌ FAIL: n parameter incorrect");
                errors = errors + 1;
            end else $display("✅ PASS: n=24 parameter correct");
            
            // Input validation - MOST CRITICAL
            if (input_a !== 32'd12345) begin
                $display("❌ CRITICAL FAIL: Input A=%0d, expected 12345", $signed(input_a));
                errors = errors + 1;
            end else $display("✅ PASS: Input A=12345 correct");
            
            if (input_b !== 32'd6789) begin
                $display("❌ CRITICAL FAIL: Input B=%0d, expected 6789", $signed(input_b));
                errors = errors + 1;
            end else $display("✅ PASS: Input B=6789 correct");
            
            // Multiplication validation
            if (mult_result_low !== 32'd83810205) begin
                $display("❌ CRITICAL FAIL: A*B=%0d, expected 83810205", $signed(mult_result_low));
                errors = errors + 1;
            end else $display("✅ PASS: Multiplication A*B=83810205 correct");
            
            if (mult_result_high !== 32'd0) begin
                $display("⚠️  WARNING: Upper 32 bits=%0d, expected 0", $signed(mult_result_high));
                warnings = warnings + 1;
            end else $display("✅ PASS: Upper 32 bits = 0 correct");
            
            // Algorithm completion validation
            if (test_counter !== 32'd5) begin
                $display("❌ FAIL: Test counter=%0d, expected 5", test_counter);
                errors = errors + 1;
            end else $display("✅ PASS: Test counter=5 algorithm completed");
            
            if (k2red_result == 32'd0) begin
                $display("⚠️  WARNING: K²RED result is 0, algorithm may be incomplete");
                warnings = warnings + 1;
            end else $display("✅ PASS: K²RED algorithm produced result=%0d", $signed(k2red_result));
            
            $display("\n📈 PERFORMANCE METRICS:");
            $display("  Total execution cycles: %0d", cyc);
            $display("  Pipeline stages: 6");
            $display("  Instructions with NOPs: 65");
            $display("  Clock frequency: 50 MHz");
            $display("  Execution time: %0d ns", cyc * 20);
            
            $display("\n🎯 DILITHIUM vs KYBER COMPARISON:");
            $display("  Kyber:     P=3329,    k=13,   m=8,  n=12");
            $display("  Dilithium: P=8380417, k=1023, m=13, n=24");
            if (p_param == 8380417 && k_param == 1023) begin
                $display("  Scale:     P is %0dx larger, k is %0dx larger", 
                         8380417/3329, 1023/13);
            end
            
            $display("\n📋 FINAL TEST SUMMARY:");
            $display("  ✅ Parameter Validation: %s", (k_param==1023 && p_param==8380417 && m_param==13 && n_param==24) ? "PASSED" : "FAILED");
            $display("  ✅ Input Validation:     %s", (input_a==12345 && input_b==6789) ? "PASSED" : "FAILED");  
            $display("  ✅ Multiplication:       %s", (mult_result_low==83810205) ? "PASSED" : "FAILED");
            $display("  ✅ Algorithm Execution:  %s", (k2red_result!=0 && test_counter==5) ? "PASSED" : "FAILED");
            $display("  📊 Total Errors: %0d", errors);
            $display("  ⚠️  Total Warnings: %0d", warnings);
            
            if (errors == 0) begin
                $display("\n🎉 SUCCESS: ALL K²RED DILITHIUM TESTS PASSED!");
                $display("✅ 6-stage pipeline synchronized correctly");
                $display("✅ Input values A=12345, B=6789 loaded properly");
                $display("✅ Multiplication 12345*6789=83810205 computed correctly");
                $display("✅ K²RED algorithm executed successfully");
                $display("✅ Test validation completed (counter=5)");
                $display("✅ Ready for CRYSTALS-Dilithium implementation");
                
                if (warnings > 0) begin
                    $display("\n⚠️  NOTE: %0d warnings detected but tests still passed", warnings);
                end
            end else begin
                $display("\n❌ FAILURE: %0d CRITICAL ERROR(S) DETECTED!", errors);
                $display("❌ Check instruction memory encoding");
                $display("❌ Verify pipeline timing and forwarding");
                $display("❌ Debug input value loading sequence");
                
                if (input_a != 12345 || input_b != 6789) begin
                    $display("\n🔧 DEBUGGING HINTS:");
                    $display("  - Input values wrong: Check LUI/ADDI instruction encoding");
                    $display("  - Verify immediate value sign extension");
                    $display("  - Check pipeline register forwarding");
                end
            end
            
            $display("\n" + "="*80);
        end
    endtask

    //---------------------------- 13. Program Termination (SYNCHRONIZED) ------
    integer program_ended;
    integer ecall_detected;
    integer ecall_cycle;
    
    initial begin
        program_ended = 0;
        ecall_detected = 0;
        ecall_cycle = 0;
    end
    
    always @(posedge clk) begin
        if (!rst && !program_ended) begin
            // Detect ECALL instruction
            if (dut.InstrD == 32'h00000073 && !ecall_detected) begin
                ecall_detected = 1;
                ecall_cycle = cyc;
                $display("\n🎯 ECALL DETECTED at cycle %0d - Dilithium algorithm complete", cyc);
                $display("📍 ECALL at PC=0x%08h (expected: 0x000000A0)", dut.PCD);
            end
            
            // Terminate after ECALL with proper 6-stage pipeline settlement
            if (ecall_detected && (cyc >= ecall_cycle + 10)) begin  // 10 cycles for 6-stage settlement
                program_ended = 1;
                $display("\n🏁 K²RED DILITHIUM TESTS COMPLETED at cycle %0d", cyc);
                repeat (3) @(posedge clk);   // Final settlement
                
                verify_dilithium_results();
                
                $fclose(trace_log);
                $display("\n🎭 SIMULATION COMPLETE - Check results above");
                $finish;
            end
            
            // UPDATED: PC range check for new instruction memory layout with extended NOPs
            if (dut.PCD > 32'h00000120) begin  // EXTENDED: Beyond ECALL at 0x110, allow more room
                program_ended = 1;
                $display("\n⚠️  PROGRAM ENDED (PC out of range) at cycle %0d", cyc);
                $display("📍 Final PC: 0x%08h (exceeded expected range 0x00000120)", dut.PCD);
                $display("🔍 This may indicate successful completion or runaway execution");
                repeat (3) @(posedge clk);
                verify_dilithium_results();
                $fclose(trace_log);
                $finish;
            end
        end
    end

    //---------------------------- 14. Safety Timeout (EXTENDED) ---------------
    initial begin
        #300000; // 300us timeout for 6-stage pipeline with NOPs
        $display("\n🚨 ERROR: Simulation timeout after 300us");
        $display("💀 Program appears to be stuck or running too long");
        $display("🔍 Final state at timeout:");
        $display("  📍 PC: 0x%08h", dut.PCD);
        $display("  📋 Current instruction: 0x%08h", dut.InstrD);
        $display("  ⏱️  Cycles executed: %0d", cyc);
        $display("  🎯 Expected completion: ~100-150 cycles");
        
        verify_dilithium_results();
        $fclose(trace_log);
        $display("\n💀 SIMULATION TERMINATED DUE TO TIMEOUT");
        $finish;
    end

    //---------------------------- 15. Early Debug (EXTENDED) ------------------
    always @(posedge clk) begin
        if (!rst && (cyc <= 75)) begin  // Extended early debug
            $display("EARLY: cyc=%0d PC=0x%08h instr=0x%08h", 
                     cyc, dut.PCD, dut.InstrD);
        end
    end

    //---------------------------- 16. Progress Indicators ----------------------
    always @(posedge clk) begin
        if (!rst && (cyc % 50 == 0) && (cyc > 0)) begin
            $display("\n⏱️  PROGRESS: Cycle %0d - Phase %0d - PC=0x%08h", 
                     cyc, test_phase, dut.PCD);
            
            // Show key register states
            if (dut.Decode.rf.regf[14] != 0 || dut.Decode.rf.regf[15] != 0) begin
                $display("📊 Key Values: A=%0d, B=%0d, A*B=%0d, Result=%0d", 
                         $signed(dut.Decode.rf.regf[14]), $signed(dut.Decode.rf.regf[15]),
                         $signed(dut.Decode.rf.regf[16]), $signed(dut.Decode.rf.regf[24]));
            end
        end
    end

    //---------------------------- 17. Critical Value Alerts (UPDATED) ----------
    always @(posedge clk) begin
        if (!rst) begin
            // Alert when key values are loaded
            if (debug_reg_write && debug_reg_addr == 5'd14 && debug_alu_result == 32'd12345) begin
                $display("\n🎯 MILESTONE: Input A=12345 loaded correctly at cycle %0d", cyc);
                $display("✅ SUCCESS: Extended NOPs fixed the A value loading!");
            end else if (debug_reg_write && debug_reg_addr == 5'd14 && debug_alu_result != 32'd12345 && debug_alu_result != 32'd0) begin
                $display("\n❌ CRITICAL: Input A=%0d (expected 12345) at cycle %0d", $signed(debug_alu_result), cyc);
                $display("🔧 Pipeline timing issue - need more NOPs or different approach");
            end
            
            if (debug_reg_write && debug_reg_addr == 5'd15 && debug_alu_result == 32'd6789) begin
                $display("🎯 MILESTONE: Input B=6789 loaded correctly at cycle %0d", cyc);
                $display("✅ SUCCESS: Extended NOPs fixed the B value loading!");
            end else if (debug_reg_write && debug_reg_addr == 5'd15 && debug_alu_result != 32'd6789 && debug_alu_result != 32'd0) begin
                $display("\n❌ CRITICAL: Input B=%0d (expected 6789) at cycle %0d", $signed(debug_alu_result), cyc);
                $display("🔧 Pipeline timing issue - check ADDI encoding");
            end
            
            if (debug_reg_write && debug_reg_addr == 5'd16 && debug_alu_result == 32'd83810205) begin
                $display("🎯 MILESTONE: Multiplication A*B=83810205 computed at cycle %0d", cyc);
                $display("✅ SUCCESS: Input values are correct and multiplication working!");
            end
            if (debug_reg_write && debug_reg_addr == 5'd24 && debug_alu_result != 32'd0) begin
                $display("🎯 MILESTONE: K²RED algorithm completed with result=%0d at cycle %0d", 
                         $signed(debug_alu_result), cyc);
            end
        end
    end

endmodule